-------------------------------------------------------------------------------
--
-- Title       : rs_trigger
-- Design      : lab_1_mks
-- Author      : maksym.popov.ki.2021@lpnu.ua
-- Company     : Lviv Polytechnic National University
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\lab_1_mks\src\Flip_Flop.vhd
-- Generated   : Mon Apr 10 20:28:56 2023
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {rs_trigger} architecture {Behavioral}}

library IEEE;
use IEEE.std_logic_1164.all;

entity rs_trigger is
	 port(
		 R : in STD_LOGIC;
		 S : in STD_LOGIC;
		 Q : out STD_LOGIC;
		 NQ : out STD_LOGIC
	     );
end rs_trigger;

--}} End of automatically maintained section

architecture Behavioral of rs_trigger is
begin

	 -- enter your statements here --

end Behavioral;
